module Input_Controller (


    
);

endmodule